// mvp Version 2.24
// cmd line +define: MIPS_SIMULATION
// cmd line +define: MIPS_VMC_DUAL_INST
// cmd line +define: MIPS_VMC_INST
// cmd line +define: M14K_NO_ERROR_GEN
// cmd line +define: M14K_NO_SHADOW_CACHE_CHECK
// cmd line +define: M14K_TRACER_NO_FDCTRACE

// Description:    m14k_clock_nogate
//       This is a replacement module for the normal toplevel clock
//       clock-gating module. Use this module for FPGA implementations.
//
//  $Id: \$
//  mips_repository_id: m14k_clock_nogate.mv, v 1.6 
//


//      	mips_start_of_legal_notice
//      	**********************************************************************
//		
//	Copyright (c) 2019 MIPS Tech, LLC, 300 Orchard City Dr., Suite 170, 
//	Campbell, CA 95008 USA.  All rights reserved.
//	This document contains information and code that is proprietary to 
//	MIPS Tech, LLC and MIPS' affiliates, as applicable, ("MIPS").  If this 
//	document is obtained pursuant to a MIPS Open license, the sole 
//	licensor under such license is MIPS Tech, LLC. This document and any 
//	information or code therein are protected by patent, copyright, 
//	trademarks and unfair competition laws, among others, and are 
//	distributed under a license restricting their use. MIPS has 
//	intellectual property rights, including patents or pending patent 
//	applications in the U.S. and in other countries, relating to the 
//	technology embodied in the product that is described in this document. 
//	Any distribution release of this document may include or be 
//	accompanied by materials developed by third parties. Any copying, 
//	reproducing, modifying or use of this information (in whole or in part) 
//	that is not expressly permitted in writing by MIPS or an authorized 
//	third party is strictly prohibited.  Any document provided in source 
//	format (i.e., in a modifiable form such as in FrameMaker or 
//	Microsoft Word format) may be subject to separate use and distribution 
//	restrictions applicable to such document. UNDER NO CIRCUMSTANCES MAY A 
//	DOCUMENT PROVIDED IN SOURCE FORMAT BE DISTRIBUTED TO A THIRD PARTY IN 
//	SOURCE FORMAT WITHOUT THE EXPRESS WRITTEN PERMISSION OF, OR LICENSED 
//	FROM, MIPS.  MIPS reserves the right to change the information or code 
//	contained in this document to improve function, design or otherwise.  
//	MIPS does not assume any liability arising out of the application or 
//	use of this information, or of any error or omission in such 
//	information. DOCUMENTATION AND CODE ARE PROVIDED "AS IS" AND ANY 
//	WARRANTIES, WHETHER EXPRESS, STATUTORY, IMPLIED OR OTHERWISE, 
//	INCLUDING BUT NOT LIMITED TO THE IMPLIED WARRANTIES OF MERCHANTABILITY, 
//	FITNESS FOR A PARTICULAR PURPOSE OR NON-INFRINGEMENT, ARE EXCLUDED, 
//	EXCEPT TO THE EXTENT THAT SUCH DISCLAIMERS ARE HELD TO BE LEGALLY 
//	INVALID IN A COMPETENT JURISDICTION. Except as expressly provided in 
//	any written license agreement from MIPS or an authorized third party, 
//	the furnishing or distribution of this document does not give recipient 
//	any license to any intellectual property rights, including any patent 
//	rights, that cover the information in this document.  
//	Products covered by, and information or code, contained this document 
//	are controlled by U.S. export control laws and may be subject to the 
//	expert or import laws in other countries. The information contained 
//	in this document shall not be exported, reexported, transferred, or 
//	released, directly or indirectly, in violation of the law of any 
//	country or international law, regulation, treaty, executive order, 
//	statute, amendments or supplements thereto. Nuclear, missile, chemical 
//	weapons, biological weapons or nuclear maritime end uses, whether 
//	direct or indirect, are strictly prohibited.  Should a conflict arise 
//	regarding the export, reexport, transfer, or release of the information 
//	contained in this document, the laws of the United States of America 
//	shall be the governing law.  
//	U.S Government Rights - Commercial software.  Government users are 
//	subject to the MIPS Tech, LLC standard license agreement and applicable 
//	provisions of the FAR and its supplements.
//	MIPS and MIPS Open are trademarks or registered trademarks of MIPS in 
//	the United States and other countries.  All other trademarks referred 
//	to herein are the property of their respective owners.  
//      
//      
//	**********************************************************************
//	mips_end_of_legal_notice
//      
////////////////////////////////////////////////////////////////////////////////

// Comments for verilint
// This is a stub module so most of the inputs are unused
//verilint 240 off  // Unused input
//verilint 528 off        // Variable set but not used

`include "m14k_const.vh"
module m14k_clock_nogate(
	gclk,
	gfclk,
	cpz_goodnight,
	SI_ClkIn,
	gscanmode,
	grfclk,
	r_gtlbclk,
	mpc_rfwrite_w,
	r_jtlb_wr,
	greset,
	jtlb_wr,
	gtlbclk);


   output 	 gclk;
   output 	 gfclk;		// Free running core clock - cannot be gated off
   input 	 cpz_goodnight;	// When Asserted, gate off the clock
   input 	 SI_ClkIn;	// Core input Clock
   input 	 gscanmode;	// When asserted, ignore cpz_goodnight and keep clock running

   output        grfclk;        // gated clock to GPRs
   output        r_gtlbclk;        // gated clock to GPRs
   input         mpc_rfwrite_w; // register write enable
   input         r_jtlb_wr;       // Write entrylo1 into the JTLB
   input	 greset;		// reset/coldreset signal
   input         jtlb_wr;       // Write entrylo1 into the JTLB
   output        gtlbclk;        // gated clock to GPRs

// BEGIN Wire declarations made by MVP
wire tracer_cg_on;
// END Wire declarations made by MVP

      
//   
   // gfclk is a buffered version of SysClk
   `M14K_CLK_BUF_CLOCK_GATE buff_fclk (	.y	(gfclk),
					.a	(SI_ClkIn)
				      );

   // gclk is also a buffered version of SysClk when no gated clocks
   `M14K_CLK_BUF_CLOCK_GATE buff_gclk (	.y	(gclk),
					.a	(SI_ClkIn)
				      );

   `M14K_CLK_BUF_CLOCK_GATE buff_gtlbclk (	.y	(gtlbclk),
					.a	(SI_ClkIn)
				      );
   `M14K_CLK_BUF_CLOCK_GATE r_buff_gtlbclk (	.y	(r_gtlbclk),
					.a	(SI_ClkIn)
				      );

    `M14K_CLK_BUF_CLOCK_GATE buff_grfclk (	.y	(grfclk),
					.a	(SI_ClkIn)
				      );

//

//verilint 599 off
//verilint 239 off
	
	assign tracer_cg_on = 1'b0;

//verilint 599 on
//verilint 239 on
//verilint 528 on        // Variable set but not used



//verilint 240 on  // Unused input

endmodule
