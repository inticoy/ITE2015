// mvp Version 2.24
// cmd line +define: MIPS_SIMULATION
// cmd line +define: MIPS_VMC_DUAL_INST
// cmd line +define: MIPS_VMC_INST
// cmd line +define: M14K_NO_ERROR_GEN
// cmd line +define: M14K_NO_SHADOW_CACHE_CHECK
// cmd line +define: M14K_TRACER_NO_FDCTRACE
//
//	Description: m14k_bistctl
//           Place-holder module for instantiation of bist controller
//
//	$Id: \$
//	mips_repository_id: m14k_bistctl.mv, v 1.1 
//

//      	mips_start_of_legal_notice
//      	**********************************************************************
//		
//	Copyright (c) 2019 MIPS Tech, LLC, 300 Orchard City Dr., Suite 170, 
//	Campbell, CA 95008 USA.  All rights reserved.
//	This document contains information and code that is proprietary to 
//	MIPS Tech, LLC and MIPS' affiliates, as applicable, ("MIPS").  If this 
//	document is obtained pursuant to a MIPS Open license, the sole 
//	licensor under such license is MIPS Tech, LLC. This document and any 
//	information or code therein are protected by patent, copyright, 
//	trademarks and unfair competition laws, among others, and are 
//	distributed under a license restricting their use. MIPS has 
//	intellectual property rights, including patents or pending patent 
//	applications in the U.S. and in other countries, relating to the 
//	technology embodied in the product that is described in this document. 
//	Any distribution release of this document may include or be 
//	accompanied by materials developed by third parties. Any copying, 
//	reproducing, modifying or use of this information (in whole or in part) 
//	that is not expressly permitted in writing by MIPS or an authorized 
//	third party is strictly prohibited.  Any document provided in source 
//	format (i.e., in a modifiable form such as in FrameMaker or 
//	Microsoft Word format) may be subject to separate use and distribution 
//	restrictions applicable to such document. UNDER NO CIRCUMSTANCES MAY A 
//	DOCUMENT PROVIDED IN SOURCE FORMAT BE DISTRIBUTED TO A THIRD PARTY IN 
//	SOURCE FORMAT WITHOUT THE EXPRESS WRITTEN PERMISSION OF, OR LICENSED 
//	FROM, MIPS.  MIPS reserves the right to change the information or code 
//	contained in this document to improve function, design or otherwise.  
//	MIPS does not assume any liability arising out of the application or 
//	use of this information, or of any error or omission in such 
//	information. DOCUMENTATION AND CODE ARE PROVIDED "AS IS" AND ANY 
//	WARRANTIES, WHETHER EXPRESS, STATUTORY, IMPLIED OR OTHERWISE, 
//	INCLUDING BUT NOT LIMITED TO THE IMPLIED WARRANTIES OF MERCHANTABILITY, 
//	FITNESS FOR A PARTICULAR PURPOSE OR NON-INFRINGEMENT, ARE EXCLUDED, 
//	EXCEPT TO THE EXTENT THAT SUCH DISCLAIMERS ARE HELD TO BE LEGALLY 
//	INVALID IN A COMPETENT JURISDICTION. Except as expressly provided in 
//	any written license agreement from MIPS or an authorized third party, 
//	the furnishing or distribution of this document does not give recipient 
//	any license to any intellectual property rights, including any patent 
//	rights, that cover the information in this document.  
//	Products covered by, and information or code, contained this document 
//	are controlled by U.S. export control laws and may be subject to the 
//	expert or import laws in other countries. The information contained 
//	in this document shall not be exported, reexported, transferred, or 
//	released, directly or indirectly, in violation of the law of any 
//	country or international law, regulation, treaty, executive order, 
//	statute, amendments or supplements thereto. Nuclear, missile, chemical 
//	weapons, biological weapons or nuclear maritime end uses, whether 
//	direct or indirect, are strictly prohibited.  Should a conflict arise 
//	regarding the export, reexport, transfer, or release of the information 
//	contained in this document, the laws of the United States of America 
//	shall be the governing law.  
//	U.S Government Rights - Commercial software.  Government users are 
//	subject to the MIPS Tech, LLC standard license agreement and applicable 
//	provisions of the FAR and its supplements.
//	MIPS and MIPS Open are trademarks or registered trademarks of MIPS in 
//	the United States and other countries.  All other trademarks referred 
//	to herein are the property of their respective owners.  
//      
//      
//	**********************************************************************
//	mips_end_of_legal_notice
//      
////////////////////////////////////////////////////////////////////////////////

// Comments for verilint...Since this is a placeholder module for bist,
//  some inputs are unused.
//verilint 240 off // Unused input

`include "m14k_const.vh"
module m14k_bistctl(
	BistIn,
	dc_bistfrom,
	ic_bistfrom,
	tcb_bistfrom,
	rf_bistfrom,
	BistOut,
	bc_dbistto,
	bc_ibistto,
	bc_tcbbistto,
	bc_rfbistto);


	/* Inputs */
	input [`M14K_TOP_BIST_IN-1:0]	BistIn;		// top-level bist input signals
	input [`M14K_DC_BIST_FROM-1:0]	dc_bistfrom;	// bist signals from dcache
	input [`M14K_IC_BIST_FROM-1:0]	ic_bistfrom;	// bist signals from icache
	input [`M14K_TCB_TRMEM_BIST_FROM-1:0]	tcb_bistfrom;	// bist signals from tcb onchip mem
	input [`M14K_RF_BIST_FROM-1:0]	rf_bistfrom;	// bist signals from generator based RF

	/* Outputs */
	output [`M14K_TOP_BIST_OUT-1:0]	BistOut;	// top-level bist output signals
	output [`M14K_DC_BIST_TO-1:0]	bc_dbistto;	// bist signals to dcache
	output [`M14K_IC_BIST_TO-1:0]	bc_ibistto;	// bist signals to icache
	output [`M14K_TCB_TRMEM_BIST_TO-1:0]	bc_tcbbistto;	// bist signals to tcb onchip mem
	output [`M14K_RF_BIST_TO-1:0]	bc_rfbistto;	// bist signals to generator based RF

// BEGIN Wire declarations made by MVP
wire [`M14K_RF_BIST_TO-1:0] /*[0:0]*/ bc_rfbistto;
wire [`M14K_DC_BIST_TO-1:0] /*[0:0]*/ bc_dbistto;
wire [`M14K_TCB_TRMEM_BIST_TO-1:0] /*[0:0]*/ bc_tcbbistto;
wire [`M14K_IC_BIST_TO-1:0] /*[0:0]*/ bc_ibistto;
wire [`M14K_TOP_BIST_OUT-1:0] /*[0:0]*/ BistOut;
// END Wire declarations made by MVP


	/* Inouts */

	// End of I/O


	/* Internal Block Wires */


	assign BistOut [`M14K_TOP_BIST_OUT-1:0] = {`M14K_TOP_BIST_OUT{1'b0}};
	assign bc_dbistto [`M14K_DC_BIST_TO-1:0] = {`M14K_DC_BIST_TO{1'b0}};
	assign bc_ibistto [`M14K_IC_BIST_TO-1:0] = {`M14K_IC_BIST_TO{1'b0}};
	assign bc_tcbbistto [`M14K_TCB_TRMEM_BIST_TO-1:0] = {`M14K_TCB_TRMEM_BIST_TO{1'b0}};
	assign bc_rfbistto [`M14K_RF_BIST_TO-1:0] = {`M14K_RF_BIST_TO{1'b0}};

//verilint 240 on // Unused input

endmodule	// m14k_bistctl
